//////////////////////////////////////////////////////////////// 
// Engineer: Evan Apinis
// 
// Module Name: instruct_mem.v
// Project Name: RV32I 
// Description: 
// 
// Instruction memory for RV32I
// 
//
// Revision 0.01 - File Created
// 
////////////////////////////////////////////////////////////////

module instruction_mem #(
  parameter MEM_SIZE = 128 // Mem size in words
)(
  input   wire        Clk_Core,
  input   wire        Rst_Core_N,
  input   wire [31:0] Program_Count,
  output  wire [31:0] Instruction
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

localparam ADDR_SIZE = $clog2(MEM_SIZE); // Parameterized address size based on mem size in words

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

reg [31:0] instr_mem [0:MEM_SIZE-1];  // Create BRAM
wire [ADDR_SIZE-1:0] 	rom_addr;	      // Read address net

integer i;

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

assign rom_addr = Program_Count[ADDR_SIZE+1:2]; // Assign effective address range
assign Instruction = instr_mem[rom_addr];       //Asynchronous read from instruct mem

initial begin
  for (i=0; i<MEM_SIZE; i=i+1) begin //Fill Instruct with 0 before writing from file
    instr_mem[i] = 32'b0;
  end
end

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////
/*
instruct_mem #(
  .DWIDTH()
  .MEM_SIZE(16384)
)
instruct_mem (
  .Clk_Core(),
  .Rst_Core_N(),
  .Program_Count(),
  .Instruction()
);
*/

endmodule